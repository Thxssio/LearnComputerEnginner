
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity p2 is
    Port ( a : in  STD_LOGIC;
           b : in  STD_LOGIC;
           c : in  STD_LOGIC;
           d : in  STD_LOGIC;
           w : out  STD_LOGIC);
end p2;

architecture Behavioral of p2 is

begin
	


end Behavioral;

